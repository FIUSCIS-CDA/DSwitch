///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: DSwitch (CLK=20)
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module testbench();
`include "../Test/Test.v"

///////////////////////////////////////////////////////////////////////////////////
// Inputs: clk, reset, D (1-bit)
reg clk, reset, D;
///////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////
// Output: Q (1-bit)
wire Q;
///////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////
// Component is CLOCKED
// Set clk period to 20 in wave
localparam CLK_PERIOD=20;
///////////////////////////////////////////////////////////////////////////////////

DSwitch mySwitch(
	.clk(clk),
	.reset(reset),
	.D(D),
        .Q(Q));


initial begin
/////////////////////////////////////////////////////////////////////////////
// Test: reset=1
$display("Testing reset: Q=0");
reset=1;  #(CLK_PERIOD/2);
verifyEqual(Q, 0);
/////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////
// Test: Falling edge
$display("Testing falling edge: Q=0");
reset=0;D=1; #(CLK_PERIOD/4);
verifyEqual(Q, 0);
/////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////////////////
// Test: Rising edge
$display("Testing rising edge: Q=D");
#(CLK_PERIOD/2);
verifyEqual(Q, D);
/////////////////////////////////////////////////////////////////////////////

$display("All tests passed.");
end

endmodule